module digito_Z (
    input A, input B, input C, input D, output oZ
);
    assign oZ = ~D;

endmodule