module digito_Y (
    input A, input B, input C, input D, output oZ
);
    not salida(oZ, D);

endmodule